----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 12/28/2023 01:06:53 PM
-- Design Name: 
-- Module Name: mux_4_to_1 - behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity mux_4_to_1 is
    port(D0,D1,D2,D3 : in std_logic_vector(7 downto 0);
         S   : in std_logic_vector(1 downto 0);
         O   : out std_logic_vector(7 downto 0));
end mux_4_to_1;

architecture behavioral of mux_4_to_1 is

begin
with S select
O <= D0 when "00",
     D1 when "01",
     D2 when "10",
     D3 when "11";
end behavioral;